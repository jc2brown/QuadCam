
library ieee;
use ieee.std_logic_1164.all;


library wifi;
use wifi.pkg_wifi.all;


entity cpt_wifi is
	port (
		i_wifi_miso : in typ_wifi_miso;
		o_wifi_mosi : out typ_wifi_mosi
	);		
end cpt_wifi;


architecture Behavioral of cpt_wifi is




begin



	

	

end Behavioral;

