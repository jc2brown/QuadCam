library ieee;
use ieee.std_logic_1164.all;

package pkg_wifi is


		
--	type typ_wifi_miso is record
--		rxd : std_logic;
--		gpio0 : std_logic;
--		gpio2 : std_logic;
--	end record;
--
--	constant init_wifi_miso : typ_wifi_miso := (
--		rxd => '1',
--		gpio0 => '0',
--		gpio2 => '0'
--	);
--
--
--	type typ_wifi_mosi is record
--		txd : std_logic;
--		rst : std_logic;	
--		ch_pd : std_logic;		
--	end record;
--
--	constant init_wifi_mosi : typ_wifi_mosi := (
--		txd => '1',
--		rst => '1',
--		ch_pd => '1'
--	);
--
--
--
--	component cpt_wifi is
--		port (
--			i_wifi_miso : in typ_wifi_miso;
--			o_wifi_mosi : out typ_wifi_mosi
--		);	
--	end component;

end pkg_wifi;

package body pkg_wifi is
end pkg_wifi;
